module pit_tben ();

reg clk=0;
reg start=0;
reg [31:0] theta=0;
reg [31:0] alpha=0;
reg [31:0] theta_setpoint=0;
reg [31:0] alpha_setpoint=0;
wire done=0;
wire [31:0] control_input=0;

parameter key_length = 512;
parameter data_length = 32;
parameter [2047:0] N2 = 508'h1778EB55F880F45868FCBBAA0E3411D3B134284D427EE14309C24941EB42E9B7A63200697FA831F9079F50C23D151877A764ACF0BE62040A94CF09BDDF23469;
parameter [15:0] N2_dash = 16'h6427;
parameter [2047:0] N_mont = 508'h138FD70691ED6093BA71A1D3DC302F7E24D692CDE4AEF2F0287E865E1FD0A1045DEB148374ED4722F556808B87B567C4D52A30E6A9B0240ECD87DF27F2F8BA5;
parameter [2047:0] N_plus_1_mont = 508'hA61394247DD8E660BC2132DD5DCFE7A8A930EBBC26C7DF710A66C272632786A2835382CAE13CEDE09C25B4B4A83599F04E7D9D7C28A5416448920E3D253BDF;
parameter [2047:0] N2_plus_2 = 508'h1778EB55F880F45868FCBBAA0E3411D3B134284D427EE14309C24941EB42E9B7A63200697FA831F9079F50C23D151877A764ACF0BE62040A94CF09BDDF2346B;
parameter [15:0] N2_plus_2_dash = 127'h27BD ;
parameter [2047:0] N = 256'h13611A1EC706880C740F5081ECE4FABD0866205F6DD4061577A9275E12695093;
parameter [15:0] N_dash = 127'h B265;
parameter [2047:0] random_seed = 508'hB1FEEFAFADBE9EFDBACD510261CCF4F17A5088BA4D402DC93BBA837CB4826C27A109463FAEFEF20662D96DA751B5E811E51EED0665E4F8FFEA89C610BD5FA8;
parameter [2047:0] lambda = 256'h33AD9AFCBD66C021357E2C0522629CA0B8D0DCD6C99331A360C85042AA8C348;
parameter [2047:0] N_inv_R_mont = 508'h14FFB8D29D6FFE75E4B10794BF40B6FD27039C9B7CB1F727884A229F5130ACB082C505AF92D33B2163C8C7DD4BDBE1DBC2381AE8446D13B6C97B7B8A916F80D;
parameter [2047:0] mu_mont = 256'hE228860E3E3B5BDC36E523B5A2B7FF2FCD227B92F62D4B7FDC1A8ED984BD474;
parameter [2047:0] k_p_theta = 1'h3;
parameter [2047:0] k_d_theta = 1'h5;
parameter [2047:0] k_alpha = 1'h7;
parameter [2047:0] neg_k_d_theta = 1'hB;
parameter [2047:0] neg_k_d_alpha = 1'hD;
parameter [2047:0] R2_mod_N2 = 508'hBDD0D1FC84A56B42D19C5A9DB797FA71960982BAB9EE33BB2485A3493B365A75012A71B635151A77167FAD41A5A2689667AFBC6EA822F61FBEEA76D6AE4476;
parameter [2047:0] R_mod_N2 = 508'hE4A4D91AE71222ABA4D2D0407E0E0D016F0A43B203C6C49F1EA2F0AF1A4C11D707C2412B8CEB9B41C0B2B81FFE30A51D72255E1D73C34120BD04B79BE7E4A3;

paillier_inverted_pendulum p_tben (
.clk(clk),
.start(start), 
.theta(theta),
.alpha(alpha),
.theta_setpoint(theta_setpoint),
.alpha_setpoint(alpha_setpoint),
.done(done), 
.control_input(control_input));


always 
#10 clk=~clk;

initial
begin 
#5; start = 1; theta = 20015;  alpha = 20017;  theta_setpoint = 210008;   alpha_setpoint = 0;
#10; start = 0; 

#89995; theta = 20004;  alpha = 20005;  theta_setpoint = 210001;   alpha_setpoint = 2;
end
endmodule