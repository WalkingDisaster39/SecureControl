module C5P(
  CLOCK_50_B3B,
  KEY,
  SW,
  LED,
  UART_TX,
  GPIO_0,
  HEX0,
  HEX1
  );


parameter cycles_per_sampling = 30000;
parameter key_length = 256;
parameter data_length = 32;
parameter [2047:0] N2 = 508'h1778EB55F880F45868FCBBAA0E3411D3B134284D427EE14309C24941EB42E9B7A63200697FA831F9079F50C23D151877A764ACF0BE62040A94CF09BDDF23469;
parameter N2_dash = 16'h6427;
parameter [2047:0] N_mont = 508'h138FD70691ED6093BA71A1D3DC302F7E24D692CDE4AEF2F0287E865E1FD0A1045DEB148374ED4722F556808B87B567C4D52A30E6A9B0240ECD87DF27F2F8BA5;
parameter [2047:0] N_plus_1_mont = 508'hA61394247DD8E660BC2132DD5DCFE7A8A930EBBC26C7DF710A66C272632786A2835382CAE13CEDE09C25B4B4A83599F04E7D9D7C28A5416448920E3D253BDF;
parameter [2047:0] N2_plus_2 = 508'h1778EB55F880F45868FCBBAA0E3411D3B134284D427EE14309C24941EB42E9B7A63200697FA831F9079F50C23D151877A764ACF0BE62040A94CF09BDDF2346B;
parameter [15:0]   N2_plus_2_dash = 16'h27BD;
parameter [2047:0] N = 256'h13611A1EC706880C740F5081ECE4FABD0866205F6DD4061577A9275E12695093;
parameter [15:0] N_dash = 16'h B265;
parameter [2047:0] random_seed = 508'hB1FEEFAFADBE9EFDBACD510261CCF4F17A5088BA4D402DC93BBA837CB4826C27A109463FAEFEF20662D96DA751B5E811E51EED0665E4F8FFEA89C610BD5FA8;
parameter [2047:0] lambda = 508'h33AD9AFCBD66C021357E2C0522629CA0B8D0DCD6C99331A360C85042AA8C348;
parameter [2047:0] N_inv_R_mont = 508'h14FFB8D29D6FFE75E4B10794BF40B6FD27039C9B7CB1F727884A229F5130ACB082C505AF92D33B2163C8C7DD4BDBE1DBC2381AE8446D13B6C97B7B8A916F80D;
parameter [2047:0] mu_mont = 256'hE228860E3E3B5BDC36E523B5A2B7FF2FCD227B92F62D4B7FDC1A8ED984BD474;
parameter [2047:0] k_p_theta = 32'hFFFFFFDF;
parameter [2047:0] k_d_theta = 32'hFFFFE00B;
parameter [2047:0] k_alpha = 32'hFFFFD623;
parameter [2047:0] neg_k_d_theta = 16'h1FF5;
parameter [2047:0] neg_k_d_alpha = 16'h27F3;
parameter [2047:0] R2_mod_N2 = 508'hBDD0D1FC84A56B42D19C5A9DB797FA71960982BAB9EE33BB2485A3493B365A75012A71B635151A77167FAD41A5A2689667AFBC6EA822F61FBEEA76D6AE4476;
parameter [2047:0] R_mod_N2 = 508'hE4A4D91AE71222ABA4D2D0407E0E0D016F0A43B203C6C49F1EA2F0AF1A4C11D707C2412B8CEB9B41C0B2B81FFE30A51D72255E1D73C34120BD04B79BE7E4A3;
parameter M_length = 512;


input CLOCK_50_B3B;
input [3:0] KEY;
input [3:0] SW;
output [3:0] LED;
output UART_TX;
inout [35:0] GPIO_0;
output [6:0] HEX0;
output [6:0] HEX1;

wire CLOCK_50_B3B;
wire [3:0] KEY;
wire [3:0] SW;
wire [3:0] LED;
wire UART_TX;
wire [35:0] GPIO_0;
wire [6:0] HEX0;
wire [6:0] HEX1;


wire clk; 
wire slow_clk;
reg [14:0] sampling_counter;
wire [14:0] speed_resized; 
wire [14:0] speed_clamped;
wire [10:0] theta_raw; 
wire [10:0] alpha_raw;
wire [data_length - 1:0] theta; 
wire [data_length - 1:0] alpha; 
wire [data_length - 1:0] control_input; 
wire [data_length - 1:0] speed_rounded; 
wire [data_length - 1:0] theta_setpoint;
wire reset_encoders; 
wire enable_motor; 
wire uart_out; 
reg start_spi; 
wire start_uart; 
wire start_paillier; 
wire done; 
reg done_reg;
wire [135:0] complex_spi;
wire [47:0] complex_uart;
wire [135:0] complex_out_spi;

paillier_inverted_pendulum paillier_inverted_pendulum (
    .clk(slow_clk),
    .start(start_paillier),
    .theta(theta),
    .alpha(alpha),
    .theta_setpoint (theta_setpoint),
    .alpha_setpoint (1024), //to_unsigned(1024, data_length),
    .done(/* open */),
    .control_input(control_input));

spi spi(
    .clk(slow_clk),
    .start(start_spi),
    .miso(GPIO_0[14]),
    .bus_in(complex_spi),
    .done(done),
    .sclk(GPIO_0[16]),
    .mosi(GPIO_0[12]),
    .ss(GPIO_0[20]),
    .bus_out(complex_out_spi));

  
uart uart(
    .clk(slow_clk),
    .start(start_uart),
    .bus_in(complex_uart),
    .done(/* open */),
    .serial_out(uart_out));


assign complex_uart = {((speed_clamped)),(alpha_raw),(theta_raw)};

assign complex_out_spi = {29'b 00000000000000000000000000000,theta_raw,13'b 0000000000000,alpha_raw,72'h 000000000000000000};

assign clk = CLOCK_50_B3B;
assign UART_TX = uart_out;

assign GPIO_0[10] = 1'b 1;
assign GPIO_0[18] = 1'b Z;
assign GPIO_0[22] = 1'b 0;

assign LED[0] = SW[0];
assign LED[1] = SW[1];
assign LED[2] = SW[2];
assign LED[3] = ~KEY[3];

assign reset_encoders =  ~KEY[3];
assign enable_motor = SW[0] == 1'b 1 && alpha_raw > 896 && alpha_raw < 1152 ? 1'b 1 : 1'b 0;

assign speed_rounded = control_input + 32'h 40;
assign speed_resized = speed_rounded [31:25];
assign speed_clamped = (speed_resized > 999) ? 14'h999 : (speed_resized < -999) ? -14'h999 : speed_resized ;

assign theta [10:0] = theta_raw;
assign alpha[10:0] = alpha_raw;
assign theta_setpoint = (SW[1] == 1'b1) ? 32'h0 : 32'hff;

assign start_paillier = done &  ~done_reg;
assign start_uart = start_spi & SW[2];
assign complex_spi = {16'h 0100,1'b 0,reset_encoders,reset_encoders,5'b 00011,96'h 000000000000000000000000,enable_motor, speed_clamped};


always @(posedge slow_clk) begin
    if((sampling_counter == (cycles_per_sampling - 1))) begin
      sampling_counter <= 0;
      start_spi <= 1'b 1;
    end
    else begin
      sampling_counter <= sampling_counter + 1;
      if((start_spi == 1'b 1)) begin
        start_spi <= 1'b 0;
      end
      done_reg <= done;
    end
  end


endmodule
